`include "cpu.svh"

module cpu
    (
        input logic clk_100M, clk_en, rst,
        input logic [31:0] r_data,
        output logic wr_en,
        output logic [31:0] mem_addr, w_data,
        // debug addr/data and instr are for showing CPU information
        // on the FPGA (only useful in synthesis)
        input logic [4:0] rdbg_addr,
        output logic [31:0] rdbg_data,
        output logic [31:0] instr,
        
        // Testing
        output logic [31:0] regA_data,
        output logic [31:0] regB_data
    );
    // The CPU interfaces with main memory which is enabled by the
    // inputs and outputs of this module (r_data, wr_en, mem_addr, w_data)
    // You should create the register file, flip flops, and logic implementing
    // a simple datapath so that instructions can be loaded from main memory,
    // executed, and the results can be inspected in the register file, or in
    // main memory (once lw and sw are supported). You should also create a
    // control FSM that controls the behavior of the datapath depending on the
    // instruction that is currently executing. You may want to split the CPU
    // into one or more submodules.
    //
    // We have provided modules for you to use inside the CPU. Please see
    // the following files:
    // reg_file.sv (register file), reg_en.sv (register with enable and reset),
    // reg_reset.sv (register with only reset), alu.sv (ALU)
    // Useful constants and opcodes are provided in cpu.svh, which is included
    // at the top of this file.
    //
    // Place the instruction machine code (generated by your assembler, or the
    // provided assembler) in asm/instr.mem and it will be automatically
    // loaded into main memory starting at address 0x00400000. Make sure the memory
    // file is imported into Vivado first (`./tcl.sh refresh`).
    
    // Testing fetching instructions
    
    // FLOW: Set next PC register
    logic PCWrite;
    logic [31:0] ALUResult; // Get ALUResult
    reg_en #(.INIT(`I_START_ADDRESS)) pc_reg (.clk(clk_100M), .rst(rst), .en(PCWrite), .d(ALUResult), .q(mem_addr));
    
    // FLOW: Get/write instruction register
    logic IRWrite; // IR write variable
    logic [31:0] IR_out; // Instructrion address
    reg_en instr_reg (.clk(clk_100M), .rst(rst), .en(IRWrite), .d(r_data), .q(IR_out));
    
    // FLOW: Mux for write register address
    logic write_addr;
    logic RegDst;
    mux_2_5bit write_addr_mux(.a(IR_out[20:16]), .b(IR_out[15:11]), .sel(RegDst), .f(write_addr));
    
    // FLOW: Register file
    logic RegWrite; // Register write variable
    logic [31:0] regA_out; 
    logic [31:0] regB_out;
    // logic [31:0] ALU_out;
    reg_file register_file (.clk(clk_100M), .wr_en(RegWrite), .r0_addr(IR_out[25:21]), 
    .r1_addr(IR_out[20:16]), .w_addr(write_addr), .w_data(ALUResult), .r0_data(regA_out), .r1_data(regB_out));
    
    // FLOW: Muxes for both ALU inputs
    logic [1:0] ALUSrcA;
    logic [1:0] ALUSrcB;
    logic [31:0] SrcA;
    logic [31:0] SrcB;
    logic [31:0] shamt;
    
    // FLOW: Zero-extend for shift amount
    assign shamt[4:0] = IR_out[10:6];
    assign shamt[31:5] = '0;
    
    // FLOW: Sign-extend for imm use
    logic [31:0] SignImm;
    assign SignImm[15:0]  = IR_out[15:0];
    assign SignImm[31:16] = IR_out[15];
    
    mux_4 mux_srcA (.a(mem_addr), .b(regA_out), .c(regB_out), .d(1'b1), .sel(ALUSrcA), .f(SrcA));
    mux_4 mux_srcB (.a(regB_out), .b(32'd4), .c(shamt), .d(SignImm), .sel(ALUSrcB), .f(SrcB));
    
    // FLOW: ALU 
    logic zero_flag;
    logic [3:0] ALUControl;
    alu alu_main (.x(SrcA), .y(SrcB), .op(ALUControl), .z(ALUResult), .zero(zero_flag));
    
    // FLOW: Register to hold ALU value
    // reg_en ALU_value (.clk(clk_100M), .rst(rst), .en(clk_en), .d(ALUResult), .q(ALU_out));
    
    // FLOW: Calculate next PC
    // logic PCSrc;
    // mux_2 mux_pcSrc (.a(ALUResult), .b(ALU_out), .sel(PCSrc), .f(PCNext));
    
    // FLOW: Declare controller
    controller cpu_controller (.rst(rst), 
        .clk(clk_100M), 
        .clk_en(clk_en),
        .opcode(IR_out[31:26]), 
        .funct(IR_out[5:0]), 
        .ALUSrcA(ALUSrcA),
        .ALUSrcB(ALUSrcB),
        .IRWrite(IRWrite),
        .PCWrite(PCWrite),
        .RegWrite(RegWrite),
        .RegDst(RegDst),
        .ALUControl(ALUControl));
    
endmodule
